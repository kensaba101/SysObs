module dpitest
(
);

    //import "DPI-C" function int getSoiValue (output int soi);
    //import "DPI-C" function void setSoiValue (output int soi, input int val); 
    //import "DPI-C" function int add (input int a, input int b);
    //export "DPI-C" function integer \$myRand;
    import "DPI-C" context function int dpic_line();

    import "DPI-C" context function logic getSoi(input logic soi); //input logic -> svLogic, output logic -> svlogic*
    export "DPI-C" function getSoiSV(input logic soi); 

    //import "DPI-C" context function void setSoi(input logic value, output logic soi);

    //initial $display("This is line %d, again, line %d\n", `__LINE__, dpic_line());


    logic testval; 



    
    initial begin
        testval = 1; 
    end

    

    function getSoiSV(input logic soi);
       /* verilator no_inline_task */
       getSoi(soi);
    endfunction


    //function setSoiSV(input logic value, output logic soi);
       /* verilator no_inline_task */
    //   setSoi(soi);
    //endfunction


endmodule