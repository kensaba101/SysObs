module fiapp
(
     clk, reset, 
